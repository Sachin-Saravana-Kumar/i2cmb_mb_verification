
    typedef enum bit [0] {
        I2C_READ = 1'b1,
        I2C_WRITE = 1'b0
    } i2c_op_t;