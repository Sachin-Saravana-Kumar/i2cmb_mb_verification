// class test_random extends ncsu_component;
//     function new();

//     endfunction
// endclass