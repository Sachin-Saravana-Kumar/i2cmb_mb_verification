    // typedef enum bit { WB_WRITE = 0 , WB_READ = 1 } wb_op_t;