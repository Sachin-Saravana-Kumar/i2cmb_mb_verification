// class test_reset_iicmb extends ncsu_component;
//     function new();
        
//     endfunction //new()
// endclass 

// class test_reg_addr_val_iicmb extends ncsu_component;
//     function new();
        
//     endfunction //new()
// endclass 

// class test_reg_permission_iicmb extends ncsu_component;
//     function new();
        
//     endfunction //new()
// endclass 

// class test_reg_alias_iicmb extends ncsu_component;
//     function new();
        
//     endfunction //new()
// endclass 
// class test_reg_def_iicmb extends ncsu_component;
//     function new();
        
//     endfunction //new()
// endclass 