// class test_i2cmb_rep_starts extends ncsu_component;
//     function new();
        
//     endfunction //new()
// endclass 

// class test_fsm_state extends ncsu_component;
//     function new();
        
//     endfunction //new()
// endclass 