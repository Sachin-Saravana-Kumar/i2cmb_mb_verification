class coverage extends ncsu_component;

endclass
